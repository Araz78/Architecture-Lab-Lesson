LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY Binary_Incrementer IS
  PORT(
    A : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    S : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    Carry_Out : OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
end Binary_Incrementer;

ARCHITECTURE structural OF Binary_Incrementer IS
SIGNAL Cout : STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL first : STD_LOGIC;
BEGIN
first <= '1';
HA_1 : entity work.Half_Adder(dataflow)
    PORT MAP(
      X => A(0),
      Y => first,
      S => S(0),
      C => Cout(0)
    );
    
HA_2 : entity work.Half_Adder(dataflow)
    PORT MAP(
      X => A(1),
      Y => Cout(0),
      S => S(1),
      C => Cout(1)
    );

HA_3 : entity work.Half_Adder(dataflow)
    PORT MAP(
      X => A(2),
      Y => Cout(1),
      S => S(2),
      C => Cout(2)
    );

HA_4 : entity work.Half_Adder(dataflow)
    PORT MAP(
      X => A(3),
      Y => Cout(2),
      S => S(3),
      C => Cout(3)
    );
Carry_Out <= Cout(3) & Cout(2) & Cout(1) & Cout(0);       
END structural;